
module nios2 (
	clk_clk);	

	input		clk_clk;
endmodule
